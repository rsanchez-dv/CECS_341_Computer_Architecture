`timescale 1ns / 1ps

module Reg2Loc(
    );


endmodule
